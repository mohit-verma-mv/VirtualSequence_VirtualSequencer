//linkedin Link 


/*

https://www.linkedin.com/pulse/difference-between-psequnecer-msequencer-uvm-raghuraj-s-bhat/

*/